
`define START_GREEN_PRINT $write("%c[1;32m",27); 
`define START_RED_PRINT $write("%c[1;31m",27);
`define START_BLUE_PRINT $write("%c[1;34m",27);
`define END_COLOR_PRINT $write("%c[0m",27);

